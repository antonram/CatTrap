// Initialize modules


// Initialize inputs and outputs
// btn will be select button

// Initialize cat




// NSL and SM
always @ (posedge Reset, posedge btn)
  

// initialize ALL variables
module CatTrap_top(
  input ClkPort
  input BtnC



);
